interface <name>_if;
    
    /*
       Define interface signals here...
    */

    
endinterface : <name>_if